module mcsassign
(

);

    reg [31:0] s;
    wire [31:0] o;
    
    assign o = s;
    
endmodule
